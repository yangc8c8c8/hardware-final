<<<<<<< HEAD
module JudgeModule(gameSTART,);
	input  gameSTART;
	output [9:0]score;
	
	`define gameIDLE 1'b0
	`define gamePLAY 1'b1
	
	always@(posedge clk)
	
	
=======
module JudgeModule(gameSTART,);
	input  gameSTART;
	output [9:0]score;
	
	`define gameIDLE 1'b0
	`define gamePLAY 1'b1
	
	always@(posedge clk)
	
	
>>>>>>> origin/master
endmodule